-------------------------------------------------------------------------------
-- Author: Bruno Albertini (balbertini@usp.br)
-- Module Name: hex2seg
-- Description:
-- VHDL module to convert from hex (4b) to 7-segment
-------------------------------------------------------------------------------

entity ascii_display is
    port (
      input: in   bit_vector(7 downto 0); -- ASCII 8 bits
      output: out bit_vector(7 downto 0)  -- ponto + abcdefg
    );
  end ascii_display;
  
  architecture comb of ascii_display is

    signal not_output : bit_vector(7 downto 0);

  begin
    output <= not not_output;
      with input select not_output <=
          "00000000" when "00100000", -- (space)
          "10000110" when "00100001", -- ! 
          "00100010" when "00100010", -- " 
          "01111110" when "00100011", -- # 
          "01101101" when "00100100", -- $ 
          "11010010" when "00100101", -- % 
          "01000110" when "00100110", -- & 
          "00100000" when "00100111", -- ' 
          "00101001" when "00101000", -- ( 
          "00001011" when "00101001", -- ) 
          "00100001" when "00101010", -- * 
          "01110000" when "00101011", -- + 
          "00010000" when "00101100", -- ,
          "01000000" when "00101101", -- - 
          "10000000" when "00101110", -- . 
          "01010010" when "00101111", -- / 
          "00111111" when "00110000", -- 0 
          "00000110" when "00110001", -- 1 
          "01011011" when "00110010", -- 2 
          "01001111" when "00110011", -- 3 
          "01100110" when "00110100", -- 4 
          "01101101" when "00110101", -- 5 
          "01111101" when "00110110", -- 6 
          "00000111" when "00110111", -- 7 
          "01111111" when "00111000", -- 8 
          "01101111" when "00111001", -- 9 
          "00001001" when "00111010", -- : 
          "00001101" when "00111011", -- ; 
          "01100001" when "00111100", -- < 
          "01001000" when "00111101", -- = 
          "01000011" when "00111110", -- > 
          "11010011" when "00111111", -- ? 
          "01011111" when "01000000", -- @ 
          "01110111" when "01000001", -- A 
          "01111100" when "01000010", -- B 
          "00111001" when "01000011", -- C 
          "01011110" when "01000100", -- D 
          "01111001" when "01000101", -- E 
          "01110001" when "01000110", -- F 
          "00111101" when "01000111", -- G 
          "01110110" when "01001000", -- H 
          "00110000" when "01001001", -- I 
          "00011110" when "01001010", -- J 
          "01110101" when "01001011", -- K 
          "00111000" when "01001100", -- L 
          "00010101" when "01001101", -- M 
          "00110111" when "01001110", -- N 
          "00111111" when "01001111", -- O 
          "01110011" when "01010000", -- P 
          "01101011" when "01010001", -- Q 
          "00110011" when "01010010", -- R 
          "01101101" when "01010011", -- S 
          "01111000" when "01010100", -- T 
          "00111110" when "01010101", -- U 
          "00111110" when "01010110", -- V 
          "00101010" when "01010111", -- W 
          "01110110" when "01011000", -- X 
          "01101110" when "01011001", -- Y 
          "01011011" when "01011010", -- Z 
          "00111001" when "01011011", -- [ 
          "01100100" when "01011100", -- \ 
          "00001111" when "01011101", -- ] 
          "00100011" when "01011110", -- ^ 
          "00001000" when "01011111", -- _ 
          "00000010" when "01100000", -- ` 
          "01011111" when "01100001", -- a 
          "01111100" when "01100010", -- b 
          "01011000" when "01100011", -- c 
          "01011110" when "01100100", -- d 
          "01111011" when "01100101", -- e 
          "01110001" when "01100110", -- f 
          "01101111" when "01100111", -- g 
          "01110100" when "01101000", -- h 
          "00010000" when "01101001", -- i 
          "00001100" when "01101010", -- j 
          "01110101" when "01101011", -- k 
          "00110000" when "01101100", -- l 
          "00010100" when "01101101", -- m 
          "01010100" when "01101110", -- n 
          "01011100" when "01101111", -- o 
          "01110011" when "01110000", -- p 
          "01100111" when "01110001", -- q 
          "01010000" when "01110010", -- r 
          "01101101" when "01110011", -- s 
          "01111000" when "01110100", -- t 
          "00011100" when "01110101", -- u 
          "00011100" when "01110110", -- v 
          "00010100" when "01110111", -- w 
          "01110110" when "01111000", -- x 
          "01101110" when "01111001", -- y 
          "01011011" when "01111010", -- z 
          "01000110" when "01111011", -- { 
          "00110000" when "01111100", -- | 
          "01110000" when "01111101", -- } 
          "00000001" when "01111110", -- ~ 
          "00000000" when "01111111", -- (del) 
          "00000000" when others;
  
  end architecture;