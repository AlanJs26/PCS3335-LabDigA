
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
 
 
ENTITY PixelGen IS
    PORT(
        RESET : IN STD_LOGIC; -- Entrada para reiniciar o estado do controlador
        F_CLOCK : IN STD_LOGIC; -- Entrada de clock (50 MHz)
        F_ON : IN STD_LOGIC; --Indica a regi�o ativa do frame
        F_ROW : IN STD_LOGIC_VECTOR(9 DOWNTO 0); -- �ndice da linha que est� sendo processada
        F_COLUMN : IN STD_LOGIC_VECTOR(10 DOWNTO 0); -- �ndice da coluna que est� sendo processada
        R_OUT : OUT STD_LOGIC; -- Componente R
        G_OUT : OUT STD_LOGIC; -- Componente G
        B_OUT : OUT STD_LOGIC -- Componente B
    );
 
END ENTITY PixelGen;
 
ARCHITECTURE arch OF PixelGen IS
SIGNAL RGBp : STD_LOGIC_VECTOR(2 DOWNTO 0); -- Valor atual do pixel
SIGNAL RGBn : STD_LOGIC_VECTOR(2 DOWNTO 0); -- �ltimo valor definido
BEGIN
 
    -- Cada componente deve ser ativada somente se o frame estiver na regi�o ativa
    R_OUT <= RGBp(2) AND F_ON;
    G_OUT <= RGBp(1) AND F_ON;
    B_OUT <= RGBp(0) AND F_ON;
        
    -- Define um novo valor RGB de acordo com �ndice da coluna
        RGBn <= "000" WHEN F_COLUMN = "0000000000" ELSE -- Preto (Coluna = 0)
                "001" WHEN F_COLUMN = "0001100100" ELSE -- Azul (Coluna = 100)
                "010" WHEN F_COLUMN = "0011001000" ELSE -- Verde (Coluna = 200)
                "011" WHEN F_COLUMN = "0100101100" ELSE -- Ciano (Coluna = 300)
                "100" WHEN F_COLUMN = "0110010000" ELSE -- Vermelho (Coluna = 400)
                "101" WHEN F_COLUMN = "0111110100" ELSE -- Magenta (Coluna = 500)
                "110" WHEN F_COLUMN = "1001011000" ELSE -- Amarelo (Coluna = 600)
                "111" WHEN F_COLUMN = "1010111100" ELSE -- Branco (Coluna = 700)
                RGBp; --�ltimo valor definido
    
    PROCESS(F_CLOCK, RESET)
    BEGIN
        IF (RESET = '0') THEN
            RGBp <= (others => '0');
        ELSIF RISING_EDGE(F_CLOCK) THEN
            RGBp <= RGBn;
        END IF;
    END PROCESS;
    
END ARCHITECTURE arch;
